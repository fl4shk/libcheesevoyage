`include "../include/misc_preprocs.svh"

class vector_add_cpkg;
endclass
