../../../../hw/gen/Gpu2dSimDut.sv