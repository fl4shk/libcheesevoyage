`ifndef MISC_PREPROCS_SVH
`define MISC_PREPROCS_SVH

`timescale 1ns/1ps
`default_nettype none

`endif		// MISC_PREPROCS_SVH
